// Testbench CSA testbench
module CSA_tb();
    reg [15:0] A, B;
    reg Cin;
    wire Cout;
    wire [15:0] Sum;
    
    CSA_design CSA(.A(A),.B(B),.Cin(Cin),.Cout(Cout),.Sum(Sum));
    
    initial begin
    $monitor("For A = %b and B = %b with Cin = %b, the Sum is %b and Cout = %b", A, B, Cin, Sum, Cout);
    
A=16'b0000000000010001; B=16'b0000010000011011; Cin = 0; #10;
A=16'b0000110011010001; B=16'b0010000011010011; Cin = 1; #10;
A=16'b0011001100110011; B=16'b0010000011010011; Cin = 0; #10;
A=16'b0100110011110011; B = 16'b0010000011010011; Cin = 0; #10;
A=16'b1000001100110011; B= 16'b1000100000110011; Cin = 1; #10;
A=16'b1100110011110011; B = 16'b0001001000001111; Cin = 0; #10;
A=16'b1111001001100111; B = 16'b1111000001110011; Cin = 0; #10;
A=16'b1111000110011011; B = 16'b1111000001110011; Cin = 1; #10;
A=16'b0000000011001100; B= 16'b0000001000001111; Cin = 0; #10;
A=16'b0000011001110001; B= 16'b0001010000011011; Cin = 1; #10;
A=16'b0011000110011011; B= 16'b0001010000011011; Cin = 0; #10;
A=16'b0110011001110011; B= 16'b0001000001110011; Cin = 0; #10;
A= 16'b1000001100110011; B=16'b1000010000011011; Cin = 1; #10;
A=16'b1100110011110011; B = 16'b0001010000011011; Cin = 0; #10;
A=16'b1111001001100111; B = 16'b1100000111110011; Cin = 0; #10;
A= 16'b1001100111110011; B = 16'b1111010000011011; Cin = 1; #10;

    end    
    initial begin
    #160;
    $finish;
    end

endmodule
